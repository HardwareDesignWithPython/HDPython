


package v_symbol_pack is 

 

end package;

package body v_symbol_pack is


end package body;
